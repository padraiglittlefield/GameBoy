module tb_control;

endmodule